// parameters

typedef 29491200 ClockFreq;
typedef 115200 BaudRate;

// derived types

typedef TDiv#(ClockFreq, BaudRate) BaudCycles;