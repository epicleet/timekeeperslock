import Keccak::*;

